interface clk_rst_intrfc;
    logic clk;
    logic rstn;
    
    //modport all_in( input clk, input rstn); //otan dhlwnw all_in tote exv san iput clk, rstn

endinterface : clk_rst_intrfc